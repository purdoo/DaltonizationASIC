library verilog;
use verilog.vl_types.all;
entity tb_encoder is
end tb_encoder;
